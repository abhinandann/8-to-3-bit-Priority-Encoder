* C:\Users\DELL\eSim-Workspace\8_3_priorityEncoder\8_3_priorityEncoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/03/22 12:25:00

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U9  Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ prioenc		
U10  I0 I1 I2 I3 I4 I5 I6 I7 Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ adc_bridge_8		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ q2 q1 q0 dac_bridge_3		
R2  q1 GND 1k		
R3  q0 GND 1k		
R1  q2 GND 1k		
v1  I0 GND pulse		
v2  I1 GND pulse		
v3  I2 GND pulse		
v4  I3 GND pulse		
v5  I4 GND pulse		
v6  I5 GND pulse		
v7  I6 GND pulse		
v8  I7 GND pulse		
U1  I0 plot_v1		
U2  I1 plot_v1		
U3  I2 plot_v1		
U4  I3 plot_v1		
U5  I4 plot_v1		
U6  I5 plot_v1		
U7  I6 plot_v1		
U8  I7 plot_v1		
U12  q0 plot_v1		
U13  q1 plot_v1		
U14  q2 plot_v1		

.end
